module system();










endmodule