module processor();










endmodule