module AHB_FIFO();












endmodule