module core();










endmodule