module operation_arm_to_std();











endmodule 