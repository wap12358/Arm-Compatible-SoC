module rom(
    clk,
    en,
    addr,
    data
);

input               clk;
input               en;
input   [31: 0]     addr;
output  [31: 0]     data;



endmodule;