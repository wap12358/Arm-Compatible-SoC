module operation_thumb_to_std();

















endmodule 