module AHB_processor();










endmodule