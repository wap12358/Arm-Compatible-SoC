module cmd_decoder_thumb(
    
);
















endmodule 